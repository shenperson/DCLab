
module pll (
	altpll_100k_clk_clk,
	altpll_12m_clk_clk,
	clk_clk,
	reset_reset_n);	

	output		altpll_100k_clk_clk;
	output		altpll_12m_clk_clk;
	input		clk_clk;
	input		reset_reset_n;
endmodule
