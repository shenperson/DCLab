module I2S(
    input clk,
    input rst,

    
);
    
endmodule